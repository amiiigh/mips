module WB_stage
(
	input	clk,
	input	rst
);
endmodule