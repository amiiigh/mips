module MEM_stage
(
	input	clk,
	input	rst
);
endmodule